LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY rom IS
	PORT(
		address : IN  std_logic_vector(4 DOWNTO 0);
		data_out : OUT std_logic_vector(18 DOWNTO 0));
END ENTITY rom;

ARCHITECTURE rom_arch OF rom IS
TYPE rom_type IS ARRAY(0 TO 31) OF std_logic_vector(18 DOWNTO 0);
	SIGNAL rom : rom_type := (
		0 => "0000010010111001100",
		1 => "0000100110010000000",
		2 => "0000000100001111000",
		3 =>"0100100110001001000",
		4 =>"0100001000001001001",
		5 =>"0010001000111001100",
		6 =>"0010011001010000100",
		7 =>"0010100010111001100",
		8 =>"0011100111000000011",
		9 =>"0011100111001001011",
		10 =>"0010110110010000000",
		11 =>"0011000101100000000",
		12 =>"0011011000110000000",
		13 =>"0011100110001001011",
		14 =>"0100000100001001001",
		15 =>"1000000000000000000",
		16 =>"0000000100000111000",
		17 =>"0100110101100000000",
		18 =>"0000001100010000000",
		19 =>"0101001100000000010",
		20 =>"0000000111000000000",
		21 =>"0000000111110010000",
		22 =>"0000001000000111000",
		23 =>"0100111001100000000",
		24 =>"0110010010111001100",
		25 =>"0110100110010000000",
		26 =>"0110110100000100000",
		27 =>"0111001011010000100",
		28 =>"0000110110101000000",
		29 =>"0111011010111001100",
		30 =>"0111100100010000000",
		31 =>"0000000110100000000"
		);
	
	BEGIN
           data_out <= rom(to_integer(unsigned(address)));

END rom_arch;

