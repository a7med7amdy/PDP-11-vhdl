LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY rom IS
	PORT(
		address : IN  std_logic_vector(4 DOWNTO 0);
		data_out : OUT std_logic_vector(17 DOWNTO 0));
END ENTITY rom;

ARCHITECTURE rom_arch OF rom IS
TYPE rom_type IS ARRAY(0 TO 31) OF std_logic_vector(17 DOWNTO 0);
	SIGNAL rom : rom_type := (
		0 => "000010010111001100",
		1 => "000100110010000000",
		2 => "000000100001111000",
		3 =>"100100110001001000",
		4 =>"100001000001001001",
		5 =>"010001000111001100",
		6 =>"010011001010000100",
		7 =>"010100010111001100",
		8 =>"011100111000000011",
		9 =>"011100111001001011",
		10 =>"010110110010000000",
		11 =>"011000101100000000",
		12 =>"011011000110000000",
		13 =>"011100110001001011",
		14 =>"100000100001001001",
		15 =>"000000000000000000",
		16 =>"000000100000111000",
		17 =>"100110101100000000",
		18 =>"000001100010000000",
		19 =>"101001100000000010",
		20 =>"000000111000000000",
		21 =>"000000111110010000",
		22 =>"000001000000111000",
		23 =>"100111001100000000",
		24 =>"110010010111001100",
		25 =>"110100110010000000",
		26 =>"110110100000100000",
		27 =>"111001011010000100",
		28 =>"000110110101000000",
		29 =>"111011010111001100",
		30 =>"111100100010000000",
		31 =>"000000110100000000"
		);
	
	BEGIN
           data_out <= rom(to_integer(unsigned(address)));

END rom_arch;

